`define RNOP 3'b000
`define RADD 3'b001
`define RSUB 3'b010
`define RMUL 3'b100